
module datapath (data, address, readM, writeM);
input data;
input address;
input readM;
input writeM;

reg data;
    always @(posedge clk) begin


    end
endmodule
