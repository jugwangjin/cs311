`timescale 1ns / 100ps

`define	NumBits	16

module ALU (A, B, FuncCode, C, OverflowFlag);
	input [`NumBits-1:0] A;
	input [`NumBits-1:0] B;
	input [3:0] FuncCode;
	output [`NumBits-1:0] C;
	output OverflowFlag;

	reg [`NumBits-1:0] C;
	reg OverflowFlag;

	// You can declare any variables as needed.
	/*
		YOUR VARIABLE DECLARATION...
	*/

	initial begin
		C = 0;
		OverflowFlag = 0;
	end   	

	// TODO: You should implement the functionality of ALU!
	// (HINT: Use 'always @(...) begin ... end')
	/*
		YOUR ALU FUNCTIONALITY IMPLEMENTATION...
	*/
	always @(A or B or FuncCode) begin
	  case (FuncCode)
	    4'b0000: 
		begin
		C = A + B;
		OverflowFlag = ((A[`NumBits-1] == 1'b1  && B[`NumBits-1] == 1'b1 && C[`NumBits-1] == 1'b0) || (A[`NumBits-1] == 1'b0 && B[`NumBits-1] == 1'b0 && C[`NumBits-1] == 1'b1)) ? 1 : 0;
		end // A + B signed addition
	    4'b0001:
		begin
		C = A - B;
		OverflowFlag = ((A[`NumBits-1] == 1'b0 && B[`NumBits-1] == 1'b1 && C[`NumBits-1] == 1'b1) || (A[`NumBits-1] == 1'b1 && B[`NumBits-1] == 1'b0 && C[`NumBits-1] == 1'b0))s ? 1 : 0;
		end // A - B signed subtraction
	    4'b0010: C = A; // A identity 
	    4'b0011: C = ~A; // ~A bitwise not
	    4'b0100: C = A & B; // A & B bitwise and
	    4'b0101: C = A | B; // A | B bitwise or
	    4'b0110: C = ~(A & B); // A nand B bitwise nand
	    4'b0111: C = ~(A | B); // A nor B bitwise nor
	    4'b1000: C = A ^ B; // A xor B bitwise xor
	    4'b1001: C = ~(A ^ B); // A nxor B bitwise xnor
	    4'b1010: C = A << 1; // A << 1 logical left shift
	    4'b1011: 
		begin
		C[`NumBits-2:0] = A[`NumBits-1:1];
		C[`NumBits-1] = 1'b0;  // A >> 1 logical right shift
		end
	    4'b1100: C = A << 1; // A <<< 1 arithmetic left shift
	    4'b1101:
		begin 
		C[`NumBits-2:0] = A[`NumBits-1:1];
		C[`NumBits-1] = C[`NumBits-2];  //A >>> 1 arithmetic right shift
		end
	    4'b1110: C = ~A + 1; // ~A + 1 2's complement
	    4'b1111: C = 0; // 0 zero
	    default: C = 0;
	  endcase
	  if (FuncCode[3:1] != 4'b000)
		begin
		OverflowFlag = 1'b0;
		end
	end
endmodule

